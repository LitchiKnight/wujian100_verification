package sim_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import yuu_common_pkg::*;
  import yuu_ahb_pkg::*;
  import yuu_int_pkg::*;
  import i2c_master_pkg::*;
  import i2c_slave_pkg::*;

  `include "sim_macro.svh"
  `include "sim_define.svh"

  `include "ral_dma.sv"
  `include "ral_wdt.sv"
  `include "ral_tim0.sv"
  `include "ral_pwm.sv"
  `include "ral_rtc.sv"
  `include "ral_usi0.sv"
  `include "top_reg_model.sv"

  `include "env_config.svh"
  `include "virtual_sequencer.svh"
  `include "env.svh"

  `include "memory_write_sequence.svh"
  `include "memory_read_sequence.svh"

  `include "wdt_int_seq.svh"
  `include "tim0_tim1_int_seq.svh"
  `include "rtc_int_seq.svh"
  `include "i2c_rx_int_seq.svh"

  `include "i2c_master_write_sequence.svh"
  `include "i2c_master_read_sequence.svh"
endpackage

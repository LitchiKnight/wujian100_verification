typedef enum int {
  ADDRESS_7BIT  = 7,
  ADDRESS_10BIT = 10
} slave_addr_mode_e;

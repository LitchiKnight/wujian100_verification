class i2c_slave_config extends uvm_object;
  `uvm_object_utils(i2c_slave_config)

  function new(string name = "i2c_slave_config");
    super.new(name);
  endfunction
endclass

// data/address width
`define ADDR_BITS            32
`define DATA_BITS            32

// base address
`define INST_SRAM_START_ADDR 32'h0000_0000
`define DATA_SRAM_START_ADDR 32'h2000_0000
`define DMA_REG_BASE_ADDR    32'h4000_0000
`define TIM0_REG_BASE_ADDR   32'h5000_0000
`define WDT_REG_BASE_ADDR    32'h5000_8000
`define PWM_REG_BASE_ADDR    32'h5001_C000
`define RTC_REG_BASE_ADDR    32'h6000_4000
`define USI0_REG_BASE_ADDR   32'h5002_8000

// memory size
`define INST_SRAM_SIZE       32'h8000
`define DATA_SRAM_SIZE       32'h3_0000

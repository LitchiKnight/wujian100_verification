interface uart_interface(
  input  rx,
  output tx
);
  logic rx;
  logic tx;
endinterface

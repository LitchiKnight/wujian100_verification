interface i2c_master_interface (input clk);
  logic scl;
  logic sda;
endinterface

typedef enum {
  INST_SRAM,
  DATA_SRAM
} memory_t;
